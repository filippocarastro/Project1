VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO rtcclock
  CLASS BLOCK ;
  FOREIGN rtcclock ;
  ORIGIN 0.000 0.000 ;
  SIZE 900.000 BY 600.000 ;
  PIN i_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.570 0.000 17.850 4.000 ;
    END
  END i_clk
  PIN i_hack
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.190 0.000 39.470 4.000 ;
    END
  END i_hack
  PIN i_wb_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.290 0.000 147.570 4.000 ;
    END
  END i_wb_addr[0]
  PIN i_wb_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.530 0.000 190.810 4.000 ;
    END
  END i_wb_addr[1]
  PIN i_wb_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.770 0.000 234.050 4.000 ;
    END
  END i_wb_addr[2]
  PIN i_wb_cyc
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.430 0.000 82.710 4.000 ;
    END
  END i_wb_cyc
  PIN i_wb_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.910 0.000 169.190 4.000 ;
    END
  END i_wb_data[0]
  PIN i_wb_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.350 0.000 428.630 4.000 ;
    END
  END i_wb_data[10]
  PIN i_wb_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.970 0.000 450.250 4.000 ;
    END
  END i_wb_data[11]
  PIN i_wb_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 471.590 0.000 471.870 4.000 ;
    END
  END i_wb_data[12]
  PIN i_wb_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 493.210 0.000 493.490 4.000 ;
    END
  END i_wb_data[13]
  PIN i_wb_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 514.830 0.000 515.110 4.000 ;
    END
  END i_wb_data[14]
  PIN i_wb_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 536.450 0.000 536.730 4.000 ;
    END
  END i_wb_data[15]
  PIN i_wb_data[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 558.070 0.000 558.350 4.000 ;
    END
  END i_wb_data[16]
  PIN i_wb_data[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.690 0.000 579.970 4.000 ;
    END
  END i_wb_data[17]
  PIN i_wb_data[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 601.310 0.000 601.590 4.000 ;
    END
  END i_wb_data[18]
  PIN i_wb_data[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 622.930 0.000 623.210 4.000 ;
    END
  END i_wb_data[19]
  PIN i_wb_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.150 0.000 212.430 4.000 ;
    END
  END i_wb_data[1]
  PIN i_wb_data[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 644.550 0.000 644.830 4.000 ;
    END
  END i_wb_data[20]
  PIN i_wb_data[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 666.170 0.000 666.450 4.000 ;
    END
  END i_wb_data[21]
  PIN i_wb_data[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 687.790 0.000 688.070 4.000 ;
    END
  END i_wb_data[22]
  PIN i_wb_data[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 709.410 0.000 709.690 4.000 ;
    END
  END i_wb_data[23]
  PIN i_wb_data[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 731.030 0.000 731.310 4.000 ;
    END
  END i_wb_data[24]
  PIN i_wb_data[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 752.650 0.000 752.930 4.000 ;
    END
  END i_wb_data[25]
  PIN i_wb_data[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 774.270 0.000 774.550 4.000 ;
    END
  END i_wb_data[26]
  PIN i_wb_data[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 795.890 0.000 796.170 4.000 ;
    END
  END i_wb_data[27]
  PIN i_wb_data[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 817.510 0.000 817.790 4.000 ;
    END
  END i_wb_data[28]
  PIN i_wb_data[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 839.130 0.000 839.410 4.000 ;
    END
  END i_wb_data[29]
  PIN i_wb_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.390 0.000 255.670 4.000 ;
    END
  END i_wb_data[2]
  PIN i_wb_data[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 860.750 0.000 861.030 4.000 ;
    END
  END i_wb_data[30]
  PIN i_wb_data[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 882.370 0.000 882.650 4.000 ;
    END
  END i_wb_data[31]
  PIN i_wb_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.010 0.000 277.290 4.000 ;
    END
  END i_wb_data[3]
  PIN i_wb_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.630 0.000 298.910 4.000 ;
    END
  END i_wb_data[4]
  PIN i_wb_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 320.250 0.000 320.530 4.000 ;
    END
  END i_wb_data[5]
  PIN i_wb_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.870 0.000 342.150 4.000 ;
    END
  END i_wb_data[6]
  PIN i_wb_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.490 0.000 363.770 4.000 ;
    END
  END i_wb_data[7]
  PIN i_wb_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 385.110 0.000 385.390 4.000 ;
    END
  END i_wb_data[8]
  PIN i_wb_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 406.730 0.000 407.010 4.000 ;
    END
  END i_wb_data[9]
  PIN i_wb_stb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.050 0.000 104.330 4.000 ;
    END
  END i_wb_stb
  PIN i_wb_we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 0.000 125.950 4.000 ;
    END
  END i_wb_we
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 596.000 26.130 600.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.250 596.000 113.530 600.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.990 596.000 122.270 600.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.730 596.000 131.010 600.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.470 596.000 139.750 600.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 596.000 148.490 600.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.950 596.000 157.230 600.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.590 596.000 34.870 600.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.330 596.000 43.610 600.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.070 596.000 52.350 600.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.810 596.000 61.090 600.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.550 596.000 69.830 600.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.290 596.000 78.570 600.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 596.000 87.310 600.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.770 596.000 96.050 600.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.510 596.000 104.790 600.000 ;
    END
  END io_oeb[9]
  PIN o_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.170 596.000 183.450 600.000 ;
    END
  END o_data[0]
  PIN o_data[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.370 596.000 445.650 600.000 ;
    END
  END o_data[10]
  PIN o_data[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 471.590 596.000 471.870 600.000 ;
    END
  END o_data[11]
  PIN o_data[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 497.810 596.000 498.090 600.000 ;
    END
  END o_data[12]
  PIN o_data[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.030 596.000 524.310 600.000 ;
    END
  END o_data[13]
  PIN o_data[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 550.250 596.000 550.530 600.000 ;
    END
  END o_data[14]
  PIN o_data[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.470 596.000 576.750 600.000 ;
    END
  END o_data[15]
  PIN o_data[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 602.690 596.000 602.970 600.000 ;
    END
  END o_data[16]
  PIN o_data[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 620.170 596.000 620.450 600.000 ;
    END
  END o_data[17]
  PIN o_data[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 637.650 596.000 637.930 600.000 ;
    END
  END o_data[18]
  PIN o_data[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 655.130 596.000 655.410 600.000 ;
    END
  END o_data[19]
  PIN o_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.390 596.000 209.670 600.000 ;
    END
  END o_data[1]
  PIN o_data[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 672.610 596.000 672.890 600.000 ;
    END
  END o_data[20]
  PIN o_data[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 690.090 596.000 690.370 600.000 ;
    END
  END o_data[21]
  PIN o_data[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 707.570 596.000 707.850 600.000 ;
    END
  END o_data[22]
  PIN o_data[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 725.050 596.000 725.330 600.000 ;
    END
  END o_data[23]
  PIN o_data[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 742.530 596.000 742.810 600.000 ;
    END
  END o_data[24]
  PIN o_data[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 760.010 596.000 760.290 600.000 ;
    END
  END o_data[25]
  PIN o_data[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 777.490 596.000 777.770 600.000 ;
    END
  END o_data[26]
  PIN o_data[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 794.970 596.000 795.250 600.000 ;
    END
  END o_data[27]
  PIN o_data[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 812.450 596.000 812.730 600.000 ;
    END
  END o_data[28]
  PIN o_data[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 829.930 596.000 830.210 600.000 ;
    END
  END o_data[29]
  PIN o_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.610 596.000 235.890 600.000 ;
    END
  END o_data[2]
  PIN o_data[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 847.410 596.000 847.690 600.000 ;
    END
  END o_data[30]
  PIN o_data[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 864.890 596.000 865.170 600.000 ;
    END
  END o_data[31]
  PIN o_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.830 596.000 262.110 600.000 ;
    END
  END o_data[3]
  PIN o_data[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.050 596.000 288.330 600.000 ;
    END
  END o_data[4]
  PIN o_data[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 314.270 596.000 314.550 600.000 ;
    END
  END o_data[5]
  PIN o_data[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.490 596.000 340.770 600.000 ;
    END
  END o_data[6]
  PIN o_data[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 366.710 596.000 366.990 600.000 ;
    END
  END o_data[7]
  PIN o_data[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.930 596.000 393.210 600.000 ;
    END
  END o_data[8]
  PIN o_data[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 419.150 596.000 419.430 600.000 ;
    END
  END o_data[9]
  PIN o_interrupt
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.690 596.000 165.970 600.000 ;
    END
  END o_interrupt
  PIN o_led[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.910 596.000 192.190 600.000 ;
    END
  END o_led[0]
  PIN o_led[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.110 596.000 454.390 600.000 ;
    END
  END o_led[10]
  PIN o_led[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 480.330 596.000 480.610 600.000 ;
    END
  END o_led[11]
  PIN o_led[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 506.550 596.000 506.830 600.000 ;
    END
  END o_led[12]
  PIN o_led[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 532.770 596.000 533.050 600.000 ;
    END
  END o_led[13]
  PIN o_led[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 558.990 596.000 559.270 600.000 ;
    END
  END o_led[14]
  PIN o_led[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 585.210 596.000 585.490 600.000 ;
    END
  END o_led[15]
  PIN o_led[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.130 596.000 218.410 600.000 ;
    END
  END o_led[1]
  PIN o_led[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.350 596.000 244.630 600.000 ;
    END
  END o_led[2]
  PIN o_led[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.570 596.000 270.850 600.000 ;
    END
  END o_led[3]
  PIN o_led[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.790 596.000 297.070 600.000 ;
    END
  END o_led[4]
  PIN o_led[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.010 596.000 323.290 600.000 ;
    END
  END o_led[5]
  PIN o_led[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 349.230 596.000 349.510 600.000 ;
    END
  END o_led[6]
  PIN o_led[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 375.450 596.000 375.730 600.000 ;
    END
  END o_led[7]
  PIN o_led[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 401.670 596.000 401.950 600.000 ;
    END
  END o_led[8]
  PIN o_led[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 427.890 596.000 428.170 600.000 ;
    END
  END o_led[9]
  PIN o_ppd
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.430 596.000 174.710 600.000 ;
    END
  END o_ppd
  PIN o_sseg[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.650 596.000 200.930 600.000 ;
    END
  END o_sseg[0]
  PIN o_sseg[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 462.850 596.000 463.130 600.000 ;
    END
  END o_sseg[10]
  PIN o_sseg[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.070 596.000 489.350 600.000 ;
    END
  END o_sseg[11]
  PIN o_sseg[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 515.290 596.000 515.570 600.000 ;
    END
  END o_sseg[12]
  PIN o_sseg[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 541.510 596.000 541.790 600.000 ;
    END
  END o_sseg[13]
  PIN o_sseg[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 567.730 596.000 568.010 600.000 ;
    END
  END o_sseg[14]
  PIN o_sseg[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 593.950 596.000 594.230 600.000 ;
    END
  END o_sseg[15]
  PIN o_sseg[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 611.430 596.000 611.710 600.000 ;
    END
  END o_sseg[16]
  PIN o_sseg[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 628.910 596.000 629.190 600.000 ;
    END
  END o_sseg[17]
  PIN o_sseg[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 646.390 596.000 646.670 600.000 ;
    END
  END o_sseg[18]
  PIN o_sseg[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 663.870 596.000 664.150 600.000 ;
    END
  END o_sseg[19]
  PIN o_sseg[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.870 596.000 227.150 600.000 ;
    END
  END o_sseg[1]
  PIN o_sseg[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 681.350 596.000 681.630 600.000 ;
    END
  END o_sseg[20]
  PIN o_sseg[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 698.830 596.000 699.110 600.000 ;
    END
  END o_sseg[21]
  PIN o_sseg[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 716.310 596.000 716.590 600.000 ;
    END
  END o_sseg[22]
  PIN o_sseg[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 733.790 596.000 734.070 600.000 ;
    END
  END o_sseg[23]
  PIN o_sseg[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 751.270 596.000 751.550 600.000 ;
    END
  END o_sseg[24]
  PIN o_sseg[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 768.750 596.000 769.030 600.000 ;
    END
  END o_sseg[25]
  PIN o_sseg[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 786.230 596.000 786.510 600.000 ;
    END
  END o_sseg[26]
  PIN o_sseg[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 803.710 596.000 803.990 600.000 ;
    END
  END o_sseg[27]
  PIN o_sseg[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 821.190 596.000 821.470 600.000 ;
    END
  END o_sseg[28]
  PIN o_sseg[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 838.670 596.000 838.950 600.000 ;
    END
  END o_sseg[29]
  PIN o_sseg[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.090 596.000 253.370 600.000 ;
    END
  END o_sseg[2]
  PIN o_sseg[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 856.150 596.000 856.430 600.000 ;
    END
  END o_sseg[30]
  PIN o_sseg[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 873.630 596.000 873.910 600.000 ;
    END
  END o_sseg[31]
  PIN o_sseg[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.310 596.000 279.590 600.000 ;
    END
  END o_sseg[3]
  PIN o_sseg[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.530 596.000 305.810 600.000 ;
    END
  END o_sseg[4]
  PIN o_sseg[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.750 596.000 332.030 600.000 ;
    END
  END o_sseg[5]
  PIN o_sseg[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.970 596.000 358.250 600.000 ;
    END
  END o_sseg[6]
  PIN o_sseg[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 384.190 596.000 384.470 600.000 ;
    END
  END o_sseg[7]
  PIN o_sseg[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 410.410 596.000 410.690 600.000 ;
    END
  END o_sseg[8]
  PIN o_sseg[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 436.630 596.000 436.910 600.000 ;
    END
  END o_sseg[9]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.810 0.000 61.090 4.000 ;
    END
  END rst
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 587.760 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 587.760 ;
    END
  END vssd1
  OBS
      LAYER nwell ;
        RECT 5.330 583.385 894.430 586.215 ;
        RECT 5.330 577.945 894.430 580.775 ;
        RECT 5.330 572.505 894.430 575.335 ;
        RECT 5.330 567.065 894.430 569.895 ;
        RECT 5.330 561.625 894.430 564.455 ;
        RECT 5.330 556.185 894.430 559.015 ;
        RECT 5.330 550.745 894.430 553.575 ;
        RECT 5.330 545.305 894.430 548.135 ;
        RECT 5.330 539.865 894.430 542.695 ;
        RECT 5.330 534.425 894.430 537.255 ;
        RECT 5.330 528.985 894.430 531.815 ;
        RECT 5.330 523.545 894.430 526.375 ;
        RECT 5.330 518.105 894.430 520.935 ;
        RECT 5.330 512.665 894.430 515.495 ;
        RECT 5.330 507.225 894.430 510.055 ;
        RECT 5.330 501.785 894.430 504.615 ;
        RECT 5.330 496.345 894.430 499.175 ;
        RECT 5.330 490.905 894.430 493.735 ;
        RECT 5.330 485.465 894.430 488.295 ;
        RECT 5.330 480.025 894.430 482.855 ;
        RECT 5.330 474.585 894.430 477.415 ;
        RECT 5.330 469.145 894.430 471.975 ;
        RECT 5.330 463.705 894.430 466.535 ;
        RECT 5.330 458.265 894.430 461.095 ;
        RECT 5.330 452.825 894.430 455.655 ;
        RECT 5.330 447.385 894.430 450.215 ;
        RECT 5.330 441.945 894.430 444.775 ;
        RECT 5.330 436.505 894.430 439.335 ;
        RECT 5.330 431.065 894.430 433.895 ;
        RECT 5.330 425.625 894.430 428.455 ;
        RECT 5.330 420.185 894.430 423.015 ;
        RECT 5.330 414.745 894.430 417.575 ;
        RECT 5.330 409.305 894.430 412.135 ;
        RECT 5.330 403.865 894.430 406.695 ;
        RECT 5.330 398.425 894.430 401.255 ;
        RECT 5.330 392.985 894.430 395.815 ;
        RECT 5.330 387.545 894.430 390.375 ;
        RECT 5.330 382.105 894.430 384.935 ;
        RECT 5.330 376.665 894.430 379.495 ;
        RECT 5.330 371.225 894.430 374.055 ;
        RECT 5.330 365.785 894.430 368.615 ;
        RECT 5.330 360.345 894.430 363.175 ;
        RECT 5.330 354.905 894.430 357.735 ;
        RECT 5.330 349.465 894.430 352.295 ;
        RECT 5.330 344.025 894.430 346.855 ;
        RECT 5.330 338.585 894.430 341.415 ;
        RECT 5.330 333.145 894.430 335.975 ;
        RECT 5.330 327.705 894.430 330.535 ;
        RECT 5.330 322.265 894.430 325.095 ;
        RECT 5.330 316.825 894.430 319.655 ;
        RECT 5.330 311.385 894.430 314.215 ;
        RECT 5.330 305.945 894.430 308.775 ;
        RECT 5.330 300.505 894.430 303.335 ;
        RECT 5.330 295.065 894.430 297.895 ;
        RECT 5.330 289.625 894.430 292.455 ;
        RECT 5.330 284.185 894.430 287.015 ;
        RECT 5.330 278.745 894.430 281.575 ;
        RECT 5.330 273.305 894.430 276.135 ;
        RECT 5.330 267.865 894.430 270.695 ;
        RECT 5.330 262.425 894.430 265.255 ;
        RECT 5.330 256.985 894.430 259.815 ;
        RECT 5.330 251.545 894.430 254.375 ;
        RECT 5.330 246.105 894.430 248.935 ;
        RECT 5.330 240.665 894.430 243.495 ;
        RECT 5.330 235.225 894.430 238.055 ;
        RECT 5.330 229.785 894.430 232.615 ;
        RECT 5.330 224.345 894.430 227.175 ;
        RECT 5.330 218.905 894.430 221.735 ;
        RECT 5.330 213.465 894.430 216.295 ;
        RECT 5.330 208.025 894.430 210.855 ;
        RECT 5.330 202.585 894.430 205.415 ;
        RECT 5.330 197.145 894.430 199.975 ;
        RECT 5.330 191.705 894.430 194.535 ;
        RECT 5.330 186.265 894.430 189.095 ;
        RECT 5.330 180.825 894.430 183.655 ;
        RECT 5.330 175.385 894.430 178.215 ;
        RECT 5.330 169.945 894.430 172.775 ;
        RECT 5.330 164.505 894.430 167.335 ;
        RECT 5.330 159.065 894.430 161.895 ;
        RECT 5.330 153.625 894.430 156.455 ;
        RECT 5.330 148.185 894.430 151.015 ;
        RECT 5.330 142.745 894.430 145.575 ;
        RECT 5.330 137.305 894.430 140.135 ;
        RECT 5.330 131.865 894.430 134.695 ;
        RECT 5.330 126.425 894.430 129.255 ;
        RECT 5.330 120.985 894.430 123.815 ;
        RECT 5.330 115.545 894.430 118.375 ;
        RECT 5.330 110.105 894.430 112.935 ;
        RECT 5.330 104.665 894.430 107.495 ;
        RECT 5.330 99.225 894.430 102.055 ;
        RECT 5.330 93.785 894.430 96.615 ;
        RECT 5.330 88.345 894.430 91.175 ;
        RECT 5.330 82.905 894.430 85.735 ;
        RECT 5.330 77.465 894.430 80.295 ;
        RECT 5.330 72.025 894.430 74.855 ;
        RECT 5.330 66.585 894.430 69.415 ;
        RECT 5.330 61.145 894.430 63.975 ;
        RECT 5.330 55.705 894.430 58.535 ;
        RECT 5.330 50.265 894.430 53.095 ;
        RECT 5.330 44.825 894.430 47.655 ;
        RECT 5.330 39.385 894.430 42.215 ;
        RECT 5.330 33.945 894.430 36.775 ;
        RECT 5.330 28.505 894.430 31.335 ;
        RECT 5.330 23.065 894.430 25.895 ;
        RECT 5.330 17.625 894.430 20.455 ;
        RECT 5.330 12.185 894.430 15.015 ;
      LAYER li1 ;
        RECT 5.520 10.795 894.240 587.605 ;
      LAYER met1 ;
        RECT 5.520 10.240 894.240 587.760 ;
      LAYER met2 ;
        RECT 17.580 595.720 25.570 596.770 ;
        RECT 26.410 595.720 34.310 596.770 ;
        RECT 35.150 595.720 43.050 596.770 ;
        RECT 43.890 595.720 51.790 596.770 ;
        RECT 52.630 595.720 60.530 596.770 ;
        RECT 61.370 595.720 69.270 596.770 ;
        RECT 70.110 595.720 78.010 596.770 ;
        RECT 78.850 595.720 86.750 596.770 ;
        RECT 87.590 595.720 95.490 596.770 ;
        RECT 96.330 595.720 104.230 596.770 ;
        RECT 105.070 595.720 112.970 596.770 ;
        RECT 113.810 595.720 121.710 596.770 ;
        RECT 122.550 595.720 130.450 596.770 ;
        RECT 131.290 595.720 139.190 596.770 ;
        RECT 140.030 595.720 147.930 596.770 ;
        RECT 148.770 595.720 156.670 596.770 ;
        RECT 157.510 595.720 165.410 596.770 ;
        RECT 166.250 595.720 174.150 596.770 ;
        RECT 174.990 595.720 182.890 596.770 ;
        RECT 183.730 595.720 191.630 596.770 ;
        RECT 192.470 595.720 200.370 596.770 ;
        RECT 201.210 595.720 209.110 596.770 ;
        RECT 209.950 595.720 217.850 596.770 ;
        RECT 218.690 595.720 226.590 596.770 ;
        RECT 227.430 595.720 235.330 596.770 ;
        RECT 236.170 595.720 244.070 596.770 ;
        RECT 244.910 595.720 252.810 596.770 ;
        RECT 253.650 595.720 261.550 596.770 ;
        RECT 262.390 595.720 270.290 596.770 ;
        RECT 271.130 595.720 279.030 596.770 ;
        RECT 279.870 595.720 287.770 596.770 ;
        RECT 288.610 595.720 296.510 596.770 ;
        RECT 297.350 595.720 305.250 596.770 ;
        RECT 306.090 595.720 313.990 596.770 ;
        RECT 314.830 595.720 322.730 596.770 ;
        RECT 323.570 595.720 331.470 596.770 ;
        RECT 332.310 595.720 340.210 596.770 ;
        RECT 341.050 595.720 348.950 596.770 ;
        RECT 349.790 595.720 357.690 596.770 ;
        RECT 358.530 595.720 366.430 596.770 ;
        RECT 367.270 595.720 375.170 596.770 ;
        RECT 376.010 595.720 383.910 596.770 ;
        RECT 384.750 595.720 392.650 596.770 ;
        RECT 393.490 595.720 401.390 596.770 ;
        RECT 402.230 595.720 410.130 596.770 ;
        RECT 410.970 595.720 418.870 596.770 ;
        RECT 419.710 595.720 427.610 596.770 ;
        RECT 428.450 595.720 436.350 596.770 ;
        RECT 437.190 595.720 445.090 596.770 ;
        RECT 445.930 595.720 453.830 596.770 ;
        RECT 454.670 595.720 462.570 596.770 ;
        RECT 463.410 595.720 471.310 596.770 ;
        RECT 472.150 595.720 480.050 596.770 ;
        RECT 480.890 595.720 488.790 596.770 ;
        RECT 489.630 595.720 497.530 596.770 ;
        RECT 498.370 595.720 506.270 596.770 ;
        RECT 507.110 595.720 515.010 596.770 ;
        RECT 515.850 595.720 523.750 596.770 ;
        RECT 524.590 595.720 532.490 596.770 ;
        RECT 533.330 595.720 541.230 596.770 ;
        RECT 542.070 595.720 549.970 596.770 ;
        RECT 550.810 595.720 558.710 596.770 ;
        RECT 559.550 595.720 567.450 596.770 ;
        RECT 568.290 595.720 576.190 596.770 ;
        RECT 577.030 595.720 584.930 596.770 ;
        RECT 585.770 595.720 593.670 596.770 ;
        RECT 594.510 595.720 602.410 596.770 ;
        RECT 603.250 595.720 611.150 596.770 ;
        RECT 611.990 595.720 619.890 596.770 ;
        RECT 620.730 595.720 628.630 596.770 ;
        RECT 629.470 595.720 637.370 596.770 ;
        RECT 638.210 595.720 646.110 596.770 ;
        RECT 646.950 595.720 654.850 596.770 ;
        RECT 655.690 595.720 663.590 596.770 ;
        RECT 664.430 595.720 672.330 596.770 ;
        RECT 673.170 595.720 681.070 596.770 ;
        RECT 681.910 595.720 689.810 596.770 ;
        RECT 690.650 595.720 698.550 596.770 ;
        RECT 699.390 595.720 707.290 596.770 ;
        RECT 708.130 595.720 716.030 596.770 ;
        RECT 716.870 595.720 724.770 596.770 ;
        RECT 725.610 595.720 733.510 596.770 ;
        RECT 734.350 595.720 742.250 596.770 ;
        RECT 743.090 595.720 750.990 596.770 ;
        RECT 751.830 595.720 759.730 596.770 ;
        RECT 760.570 595.720 768.470 596.770 ;
        RECT 769.310 595.720 777.210 596.770 ;
        RECT 778.050 595.720 785.950 596.770 ;
        RECT 786.790 595.720 794.690 596.770 ;
        RECT 795.530 595.720 803.430 596.770 ;
        RECT 804.270 595.720 812.170 596.770 ;
        RECT 813.010 595.720 820.910 596.770 ;
        RECT 821.750 595.720 829.650 596.770 ;
        RECT 830.490 595.720 838.390 596.770 ;
        RECT 839.230 595.720 847.130 596.770 ;
        RECT 847.970 595.720 855.870 596.770 ;
        RECT 856.710 595.720 864.610 596.770 ;
        RECT 865.450 595.720 873.350 596.770 ;
        RECT 874.190 595.720 884.480 596.770 ;
        RECT 17.580 4.280 884.480 595.720 ;
        RECT 18.130 3.670 38.910 4.280 ;
        RECT 39.750 3.670 60.530 4.280 ;
        RECT 61.370 3.670 82.150 4.280 ;
        RECT 82.990 3.670 103.770 4.280 ;
        RECT 104.610 3.670 125.390 4.280 ;
        RECT 126.230 3.670 147.010 4.280 ;
        RECT 147.850 3.670 168.630 4.280 ;
        RECT 169.470 3.670 190.250 4.280 ;
        RECT 191.090 3.670 211.870 4.280 ;
        RECT 212.710 3.670 233.490 4.280 ;
        RECT 234.330 3.670 255.110 4.280 ;
        RECT 255.950 3.670 276.730 4.280 ;
        RECT 277.570 3.670 298.350 4.280 ;
        RECT 299.190 3.670 319.970 4.280 ;
        RECT 320.810 3.670 341.590 4.280 ;
        RECT 342.430 3.670 363.210 4.280 ;
        RECT 364.050 3.670 384.830 4.280 ;
        RECT 385.670 3.670 406.450 4.280 ;
        RECT 407.290 3.670 428.070 4.280 ;
        RECT 428.910 3.670 449.690 4.280 ;
        RECT 450.530 3.670 471.310 4.280 ;
        RECT 472.150 3.670 492.930 4.280 ;
        RECT 493.770 3.670 514.550 4.280 ;
        RECT 515.390 3.670 536.170 4.280 ;
        RECT 537.010 3.670 557.790 4.280 ;
        RECT 558.630 3.670 579.410 4.280 ;
        RECT 580.250 3.670 601.030 4.280 ;
        RECT 601.870 3.670 622.650 4.280 ;
        RECT 623.490 3.670 644.270 4.280 ;
        RECT 645.110 3.670 665.890 4.280 ;
        RECT 666.730 3.670 687.510 4.280 ;
        RECT 688.350 3.670 709.130 4.280 ;
        RECT 709.970 3.670 730.750 4.280 ;
        RECT 731.590 3.670 752.370 4.280 ;
        RECT 753.210 3.670 773.990 4.280 ;
        RECT 774.830 3.670 795.610 4.280 ;
        RECT 796.450 3.670 817.230 4.280 ;
        RECT 818.070 3.670 838.850 4.280 ;
        RECT 839.690 3.670 860.470 4.280 ;
        RECT 861.310 3.670 882.090 4.280 ;
        RECT 882.930 3.670 884.480 4.280 ;
      LAYER met3 ;
        RECT 21.050 10.715 867.430 587.685 ;
      LAYER met4 ;
        RECT 371.975 332.695 404.640 534.305 ;
        RECT 407.040 332.695 481.440 534.305 ;
        RECT 483.840 332.695 558.240 534.305 ;
        RECT 560.640 332.695 575.625 534.305 ;
  END
END rtcclock
END LIBRARY

